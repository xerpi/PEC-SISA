-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Fri Mar 18 16:44:29 2016

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY SM1 IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clk : IN STD_LOGIC;
        WR : IN STD_LOGIC := '0';
        byte_m : IN STD_LOGIC := '0';
        lsb : IN STD_LOGIC := '0';
        cont : IN STD_LOGIC_VECTOR(2 DOWNTO 0) := "000";
        SRAM_UB_N : OUT STD_LOGIC;
        SRAM_LB_N : OUT STD_LOGIC;
        SRAM_CE_N : OUT STD_LOGIC;
        SRAM_OE_N : OUT STD_LOGIC;
        SRAM_WE_N : OUT STD_LOGIC
    );
END SM1;

ARCHITECTURE BEHAVIOR OF SM1 IS
    TYPE type_fstate IS (READ,WRITEW,WRITEB_0,WRITEB_1);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clk,reg_fstate)
    BEGIN
        IF (clk='1' AND clk'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,WR,byte_m,lsb,cont)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= READ;
            SRAM_UB_N <= '0';
            SRAM_LB_N <= '0';
            SRAM_CE_N <= '0';
            SRAM_OE_N <= '0';
            SRAM_WE_N <= '0';
        ELSE
            SRAM_UB_N <= '0';
            SRAM_LB_N <= '0';
            SRAM_CE_N <= '0';
            SRAM_OE_N <= '0';
            SRAM_WE_N <= '0';
            CASE fstate IS
                WHEN READ =>
                    IF (NOT((WR = '1'))) THEN
                        reg_fstate <= READ;
                    ELSIF ((((WR = '1') AND NOT((byte_m = '1'))) AND (cont(2 DOWNTO 0) = "000"))) THEN
                        reg_fstate <= WRITEW;
                    ELSIF (((((WR = '1') AND (byte_m = '1')) AND NOT((lsb = '1'))) AND (cont(2 DOWNTO 0) = "000"))) THEN
                        reg_fstate <= WRITEB_0;
                    ELSIF (((((WR = '1') AND (byte_m = '1')) AND (lsb = '1')) AND (cont(2 DOWNTO 0) = "000"))) THEN
                        reg_fstate <= WRITEB_1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= READ;
                    END IF;

                    SRAM_CE_N <= '0';

                    SRAM_UB_N <= '0';

                    SRAM_WE_N <= '1';

                    SRAM_LB_N <= '0';

                    SRAM_OE_N <= '0';
                WHEN WRITEW =>
                    reg_fstate <= READ;

                    SRAM_CE_N <= '0';

                    SRAM_UB_N <= '0';

                    SRAM_WE_N <= '0';

                    SRAM_LB_N <= '0';

                    SRAM_OE_N <= '0';
                WHEN WRITEB_0 =>
                    reg_fstate <= READ;

                    SRAM_CE_N <= '0';

                    SRAM_UB_N <= '1';

                    SRAM_WE_N <= '0';

                    SRAM_LB_N <= '0';

                    SRAM_OE_N <= '0';
                WHEN WRITEB_1 =>
                    reg_fstate <= READ;

                    SRAM_CE_N <= '0';

                    SRAM_UB_N <= '0';

                    SRAM_WE_N <= '0';

                    SRAM_LB_N <= '1';

                    SRAM_OE_N <= '0';
                WHEN OTHERS => 
                    SRAM_UB_N <= 'X';
                    SRAM_LB_N <= 'X';
                    SRAM_CE_N <= 'X';
                    SRAM_OE_N <= 'X';
                    SRAM_WE_N <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
